The purpose of this dummy file is to create this directory.